library verilog;
use verilog.vl_types.all;
entity maiorQue_vlg_check_tst is
    port(
        s               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end maiorQue_vlg_check_tst;
