library verilog;
use verilog.vl_types.all;
entity inversor is
    port(
        x1              : in     vl_logic;
        Y               : out    vl_logic
    );
end inversor;
