library verilog;
use verilog.vl_types.all;
entity maiorQue_vlg_vec_tst is
end maiorQue_vlg_vec_tst;
