library verilog;
use verilog.vl_types.all;
entity Calculadora_vlg_vec_tst is
end Calculadora_vlg_vec_tst;
