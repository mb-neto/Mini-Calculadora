library verilog;
use verilog.vl_types.all;
entity inversor_vlg_sample_tst is
    port(
        x1              : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end inversor_vlg_sample_tst;
