library verilog;
use verilog.vl_types.all;
entity Subtrador_vlg_vec_tst is
end Subtrador_vlg_vec_tst;
